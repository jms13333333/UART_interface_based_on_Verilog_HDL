`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/01/27 16:04:34
// Design Name: 
// Module Name: UART_TX
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module UART_TX(
    input wire clk, 
    input wire resetn, 
    output wire uart_txd,
    output wire uart_tx_busy,
    input wire uart_tx_en, 
    input wire [7:0] uart_tx_data  
    );
    parameter BIT_RATE=9600; // bits / sec
    localparam BIT_P=1_000_000_000 * 1/BIT_RATE;
    parameter CLK_HZ=50_000_000;
    localparam CLK_P=1_000_000_000 * 1/CLK_HZ;
    parameter STOP_BITS=1;
    localparam CYCLES_PER_BIT=BIT_P / CLK_P;
    localparam COUNT_REG_LEN=1+$clog2(CYCLES_PER_BIT);
    reg txd_reg;
    reg [7:0] data_to_send;
    reg [COUNT_REG_LEN-1:0] cycle_counter;
    reg [3:0] bit_counter;
    reg [2:0] fsm_state;
    reg [2:0] n_fsm_state;
    
    localparam FSM_IDLE = 0;
    localparam FSM_START= 1;
    localparam FSM_SEND = 2;
    localparam FSM_STOP = 3;
    
    assign uart_tx_busy = fsm_state != FSM_IDLE;
    assign uart_txd     = txd_reg;
    
    wire next_bit     = cycle_counter == CYCLES_PER_BIT;
    wire payload_done = bit_counter   == 8  ;
    wire stop_done    = bit_counter   == STOP_BITS && fsm_state == FSM_STOP;
    // Handle picking the next state.
    always @(*) begin : p_n_fsm_state
        case(fsm_state)
            FSM_IDLE : n_fsm_state = uart_tx_en   ? FSM_START: FSM_IDLE ;
            FSM_START: n_fsm_state = next_bit     ? FSM_SEND : FSM_START;
            FSM_SEND : n_fsm_state = payload_done ? FSM_STOP : FSM_SEND ;
            FSM_STOP : n_fsm_state = stop_done    ? FSM_IDLE : FSM_STOP ;
            default  : n_fsm_state = FSM_IDLE;
        endcase
    end
    
    integer i = 0;
    always @(posedge clk) begin : p_data_to_send
        if(!resetn) begin
            data_to_send <= {8{1'b0}};
        end else if(fsm_state == FSM_IDLE && uart_tx_en) begin
            data_to_send <= uart_tx_data;
        end else if(fsm_state       == FSM_SEND       && next_bit ) begin
            for ( i = 6; i >= 0; i = i - 1) begin
                data_to_send[i] <= data_to_send[i+1];
            end
        end
    end
    
    always @(posedge clk) begin : p_bit_counter
        if(!resetn) begin
            bit_counter <= 4'b0;
        end else if(fsm_state != FSM_SEND && fsm_state != FSM_STOP) begin
            bit_counter <= {COUNT_REG_LEN{1'b0}};
        end else if(fsm_state == FSM_SEND && n_fsm_state == FSM_STOP) begin
            bit_counter <= {COUNT_REG_LEN{1'b0}};
        end else if(fsm_state == FSM_STOP&& next_bit) begin
            bit_counter <= bit_counter + 1'b1;
        end else if(fsm_state == FSM_SEND && next_bit) begin
            bit_counter <= bit_counter + 1'b1;
        end
    end
    
    always @(posedge clk) begin : p_cycle_counter
        if(!resetn) begin
            cycle_counter <= {COUNT_REG_LEN{1'b0}};
        end else if(next_bit) begin
            cycle_counter <= {COUNT_REG_LEN{1'b0}};
        end else if(fsm_state == FSM_START || 
                    fsm_state == FSM_SEND  || 
                    fsm_state == FSM_STOP   ) begin
            cycle_counter <= cycle_counter + 1'b1;
        end
    end
    
    always @(posedge clk) begin : p_fsm_state
        if(!resetn) begin
            fsm_state <= FSM_IDLE;
        end else begin
            fsm_state <= n_fsm_state;
        end
    end
    
    // Responsible for updating the internal value of the txd_reg.
    always @(posedge clk) begin : p_txd_reg
        if(!resetn) begin
            txd_reg <= 1'b1;
        end else if(fsm_state == FSM_IDLE) begin
            txd_reg <= 1'b1;
        end else if(fsm_state == FSM_START) begin
            txd_reg <= 1'b0;
        end else if(fsm_state == FSM_SEND) begin
            txd_reg <= data_to_send[0];
        end else if(fsm_state == FSM_STOP) begin
            txd_reg <= 1'b1;
        end
    end
endmodule
