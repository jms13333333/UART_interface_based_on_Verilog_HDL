`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/01/27 16:34:25
// Design Name: 
// Module Name: UART_TOP
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module UART_TOP(
    input clk     , // Top level system clock input.
    input sw_0    , // Slide switches.
    input sw_1    , // Slide switches.
    input wire uart_rxd, // UART Recieve pin.
    output wire uart_txd, // UART transmit pin.
    output wire [7:0] led
    );
    parameter CLK_HZ = 50000000;
    parameter BIT_RATE =   9600;
    parameter PAYLOAD_BITS = 8;
    
    wire [PAYLOAD_BITS-1:0]  uart_rx_data;
    wire uart_rx_valid;
    wire uart_rx_break;
    wire uart_tx_busy;
    wire [PAYLOAD_BITS-1:0]  uart_tx_data;
    wire uart_tx_en;
    
    reg  [PAYLOAD_BITS-1:0]  led_reg;
    assign led = led_reg;
    assign uart_tx_data = uart_rx_data;
    assign uart_tx_en   = uart_rx_valid;
    always @(posedge clk) begin
        if(!sw_0) begin
            led_reg <= 8'hF0;
        end else if(uart_rx_valid) begin
            led_reg <= uart_rx_data[7:0];
        end
    end
    
    UART_RX #(
        .BIT_RATE(BIT_RATE),
        .CLK_HZ  (CLK_HZ  )
    ) i_uart_rx(
        .clk          (clk          ), // Top level system clock input.
        .resetn       (sw_0         ), // Asynchronous active low reset.
        .uart_rxd     (uart_rxd     ), // UART Recieve pin.
        .uart_rx_en   (1'b1         ), // Recieve enable
        .uart_rx_break(uart_rx_break), // Did we get a BREAK message?
        .uart_rx_valid(uart_rx_valid), // Valid data recieved and available.
        .uart_rx_data (uart_rx_data )  // The recieved data.
    );
    UART_TX #(
        .BIT_RATE(BIT_RATE),
        .CLK_HZ  (CLK_HZ  )
        ) i_uart_tx(
        .clk          (clk          ),
        .resetn       (sw_0         ),
        .uart_txd     (uart_txd     ),
        .uart_tx_en   (uart_tx_en   ),
        .uart_tx_busy (uart_tx_busy ),
        .uart_tx_data (uart_tx_data ) 
    );
endmodule